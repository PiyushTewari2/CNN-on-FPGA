`timescale 1ns / 1ps

module conv_core_product_controller(

    );
endmodule
