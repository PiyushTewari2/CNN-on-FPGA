`timescale 1ns / 1ps

module con_core_top(

    );
endmodule
