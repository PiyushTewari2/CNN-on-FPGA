`timescale 1ns / 1ps

module conv_core_accumulator(

    );
endmodule
